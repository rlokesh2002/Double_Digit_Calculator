CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1534 795
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 1 2 1
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
73
9 2-In NOR~
219 800 870 0 3 22
0 3 4 55
0
0 0 624 782
6 74LS02
-21 -24 21 -16
3 U1A
31 -10 52 -2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 3 2 1 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 1 17 0
1 U
3557 0 0
2
44808.7 0
0
9 Inverter~
13 123 625 0 2 22
0 15 13
0
0 0 624 602
6 74LS04
-21 -19 21 -11
3 U4E
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 4 0
1 U
7246 0 0
2
44808.7 0
0
9 Inverter~
13 93 665 0 2 22
0 16 14
0
0 0 624 602
6 74LS04
-21 -19 21 -11
3 U4D
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 4 0
1 U
3916 0 0
2
44808.7 0
0
6 74LS83
105 1197 2280 0 14 29
0 2 2 7 7 31 30 29 27 2
18 19 20 21 176
0
0 0 13040 782
7 74LS83A
-24 -60 25 -52
3 U51
56 -2 77 6
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 512 1 0 0 0
1 U
614 0 0
2
44808.7 1
0
6 74LS85
106 1123 2179 0 14 29
0 2 28 2 2 31 30 29 27 177
28 178 7 179 180
0
0 0 5104 782
6 74LS85
48 3 90 11
3 U52
58 -7 79 1
0
15 DVCC=16;DGND=8;
136 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 13 12 10 1 14 11 9 2
3 4 7 6 5 15 13 12 10 1
14 11 9 2 3 4 7 6 5 0
65 0 0 512 0 0 0 0
1 U
8494 0 0
2
44808.7 0
0
6 74LS85
106 1123 1930 0 14 29
0 2 28 2 2 2 34 33 32 181
28 182 8 183 184
0
0 0 5104 782
6 74LS85
48 3 90 11
3 U49
58 -7 79 1
0
15 DVCC=16;DGND=8;
136 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 13 12 10 1 14 11 9 2
3 4 7 6 5 15 13 12 10 1
14 11 9 2 3 4 7 6 5 0
65 0 0 512 0 0 0 0
1 U
774 0 0
2
44808.7 1
0
6 74LS83
105 1197 2031 0 14 29
0 2 2 8 8 2 34 33 32 2
185 31 30 29 186
0
0 0 13040 782
7 74LS83A
-24 -60 25 -52
3 U50
56 -2 77 6
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 512 1 0 0 0
1 U
715 0 0
2
44808.7 0
0
6 74LS85
106 785 2139 0 14 29
0 2 28 2 2 38 37 36 35 187
28 188 9 189 190
0
0 0 5104 782
6 74LS85
48 3 90 11
3 U48
58 -7 79 1
0
15 DVCC=16;DGND=8;
136 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 13 12 10 1 14 11 9 2
3 4 7 6 5 15 13 12 10 1
14 11 9 2 3 4 7 6 5 0
65 0 0 512 0 0 0 0
1 U
3281 0 0
2
44808.7 1
0
6 74LS83
105 859 2240 0 14 29
0 2 2 9 9 38 37 36 35 2
22 23 24 25 191
0
0 0 13040 782
7 74LS83A
-24 -60 25 -52
3 U47
56 -2 77 6
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 512 1 0 0 0
1 U
3593 0 0
2
44808.7 0
0
6 74LS83
105 859 1995 0 14 29
0 2 2 10 10 42 41 40 39 2
27 38 37 36 192
0
0 0 13040 782
7 74LS83A
-24 -60 25 -52
3 U46
56 -2 77 6
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 512 1 0 0 0
1 U
7233 0 0
2
44808.7 1
0
6 74LS85
106 785 1894 0 14 29
0 2 28 2 2 42 41 40 39 193
28 194 10 195 196
0
0 0 5104 782
6 74LS85
48 3 90 11
3 U45
58 -7 79 1
0
15 DVCC=16;DGND=8;
136 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 13 12 10 1 14 11 9 2
3 4 7 6 5 15 13 12 10 1
14 11 9 2 3 4 7 6 5 0
65 0 0 512 0 0 0 0
1 U
3410 0 0
2
44808.7 0
0
6 74LS85
106 785 1648 0 14 29
0 2 28 2 2 46 45 44 43 197
28 198 11 199 200
0
0 0 5104 782
6 74LS85
48 3 90 11
3 U44
58 -7 79 1
0
15 DVCC=16;DGND=8;
136 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 13 12 10 1 14 11 9 2
3 4 7 6 5 15 13 12 10 1
14 11 9 2 3 4 7 6 5 0
65 0 0 512 0 0 0 0
1 U
3616 0 0
2
44808.7 1
0
6 74LS83
105 859 1749 0 14 29
0 2 2 11 11 46 45 44 43 2
32 42 41 40 201
0
0 0 13040 782
7 74LS83A
-24 -60 25 -52
3 U43
56 -2 77 6
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 512 1 0 0 0
1 U
5202 0 0
2
44808.7 0
0
6 74LS83
105 859 1502 0 14 29
0 2 2 12 12 50 49 48 47 2
33 46 45 44 202
0
0 0 13040 782
7 74LS83A
-24 -60 25 -52
3 U42
56 -2 77 6
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 512 1 0 0 0
1 U
9145 0 0
2
44808.7 1
0
6 74LS85
106 785 1401 0 14 29
0 2 28 2 2 50 49 48 47 203
28 204 12 205 206
0
0 0 5104 782
6 74LS85
48 3 90 11
3 U41
58 -7 79 1
0
15 DVCC=16;DGND=8;
136 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 13 12 10 1 14 11 9 2
3 4 7 6 5 15 13 12 10 1
14 11 9 2 3 4 7 6 5 0
65 0 0 512 0 0 0 0
1 U
9815 0 0
2
44808.7 0
0
2 +V
167 708 961 0 1 3
0 28
0
0 0 54256 0
2 5V
-8 -22 6 -14
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
4766 0 0
2
44808.7 0
0
7 Ground~
168 752 944 0 1 3
0 2
0
0 0 53360 180
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
8325 0 0
2
44808.7 0
0
6 74LS85
106 785 1160 0 14 29
0 2 28 2 2 2 52 53 54 207
28 208 51 209 210
0
0 0 5104 782
6 74LS85
48 3 90 11
3 U39
58 -7 79 1
0
15 DVCC=16;DGND=8;
136 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 13 12 10 1 14 11 9 2
3 4 7 6 5 15 13 12 10 1
14 11 9 2 3 4 7 6 5 0
65 0 0 512 0 0 0 0
1 U
7196 0 0
2
44808.7 1
0
6 74LS83
105 859 1253 0 14 29
0 2 2 51 51 2 52 53 54 2
34 50 49 48 211
0
0 0 13040 782
7 74LS83A
-24 -60 25 -52
3 U40
56 -2 77 6
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 512 1 0 0 0
1 U
3567 0 0
2
44808.7 0
0
9 2-In AND~
219 804 729 0 3 22
0 3 4 17
0
0 0 624 782
6 74LS08
-21 -24 21 -16
4 U38A
17 -4 45 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 16 0
1 U
5877 0 0
2
44808.7 0
0
7 Ground~
168 686 758 0 1 3
0 2
0
0 0 53360 180
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
4785 0 0
2
44808.7 0
0
10 3-In NAND~
219 1405 199 0 4 22
0 126 140 139 125
0
0 0 624 512
6 74LS10
-21 -28 21 -20
4 U37A
-11 -25 17 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 1 15 0
1 U
3822 0 0
2
44808.7 0
0
9 Inverter~
13 880 693 0 2 22
0 64 4
0
0 0 624 180
6 74LS04
-21 -19 21 -11
3 U4C
-5 -20 16 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 4 0
1 U
7640 0 0
2
44808.6 0
0
6 74LS83
105 877 1074 0 14 29
0 2 2 2 2 55 56 57 58 59
52 53 54 47 212
0
0 0 13040 782
7 74LS83A
-24 -60 25 -52
3 U36
56 -2 77 6
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 512 1 0 0 0
1 U
9221 0 0
2
44808.6 0
0
9 2-In XOR~
219 1073 1029 0 3 22
0 78 17 61
0
0 0 624 270
6 74LS86
-21 -24 21 -16
4 U33A
-10 -4 18 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 1 14 0
1 U
6484 0 0
2
44808.6 3
0
9 2-In XOR~
219 988 1027 0 3 22
0 76 17 63
0
0 0 624 270
6 74LS86
-21 -24 21 -16
4 U24A
-11 -3 17 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 1 8 0
1 U
3689 0 0
2
44808.6 2
0
9 2-In XOR~
219 1030 1028 0 3 22
0 77 17 62
0
0 0 624 270
6 74LS86
-21 -24 21 -16
4 U21A
-11 -1 17 7
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 1 7 0
1 U
3952 0 0
2
44808.6 1
0
9 2-In XOR~
219 1115 1029 0 3 22
0 79 17 60
0
0 0 624 270
6 74LS86
-21 -24 21 -16
4 U10A
-12 -3 16 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 1 5 0
1 U
3631 0 0
2
44808.6 0
0
9 2-In XOR~
219 935 854 0 3 22
0 75 17 58
0
0 0 624 270
6 74LS86
-21 -24 21 -16
4 U22B
-12 -3 16 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 2 12 0
1 U
9359 0 0
2
44808.6 3
0
9 2-In XOR~
219 850 853 0 3 22
0 73 17 56
0
0 0 624 270
6 74LS86
-21 -24 21 -16
4 U22C
-11 -1 17 7
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 3 12 0
1 U
5584 0 0
2
44808.6 2
0
9 2-In XOR~
219 893 854 0 3 22
0 74 17 57
0
0 0 624 270
6 74LS86
-21 -24 21 -16
3 U7A
-7 -4 14 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 1 3 0
1 U
4973 0 0
2
44808.6 0
0
6 74LS83
105 1046 1144 0 14 29
0 63 62 61 60 2 2 2 2 17
43 39 35 26 59
0
0 0 13040 782
7 74LS83A
-24 -60 25 -52
2 U8
57 -2 71 6
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 0 1 0 0 0
1 U
3239 0 0
2
44808.6 0
0
6 74LS83
105 1002 795 0 14 29
0 2 80 81 82 84 85 86 87 83
64 73 74 75 213
0
0 0 13040 512
7 74LS83A
-24 -60 25 -52
2 U5
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 512 1 0 0 0
1 U
4244 0 0
2
44808.6 0
0
6 74LS83
105 1170 950 0 14 29
0 88 89 90 91 92 93 94 95 3
76 77 78 79 83
0
0 0 13040 512
7 74LS83A
-24 -60 25 -52
2 U3
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 0 1 0 0 0
1 U
3391 0 0
2
44808.6 0
0
9 2-In XOR~
219 1076 641 0 3 22
0 3 100 82
0
0 0 624 270
6 74LS86
-21 -24 21 -16
4 U18A
-12 -2 16 6
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 1 2 0
1 U
4243 0 0
2
44808.6 3
0
9 2-In XOR~
219 991 640 0 3 22
0 3 102 80
0
0 0 624 270
6 74LS86
-21 -24 21 -16
4 U20A
-11 -1 17 7
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 1 10 0
1 U
3907 0 0
2
44808.6 2
0
9 2-In XOR~
219 1034 641 0 3 22
0 3 101 81
0
0 0 624 270
6 74LS86
-21 -24 21 -16
4 U19A
-10 -4 18 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 1 9 0
1 U
728 0 0
2
44808.6 0
0
9 2-In XOR~
219 1212 711 0 3 22
0 3 97 90
0
0 0 624 270
6 74LS86
-21 -24 21 -16
4 U15B
-10 -4 18 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 2 11 0
1 U
3585 0 0
2
44808.6 3
0
9 2-In XOR~
219 1169 710 0 3 22
0 3 98 89
0
0 0 624 270
6 74LS86
-21 -24 21 -16
4 U15C
-11 -1 17 7
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 3 11 0
1 U
3565 0 0
2
44808.6 2
0
9 2-In XOR~
219 1127 709 0 3 22
0 3 99 88
0
0 0 624 270
6 74LS86
-21 -24 21 -16
4 U15A
-11 -3 17 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 1 11 0
1 U
3966 0 0
2
44808.6 1
0
9 2-In XOR~
219 1254 711 0 3 22
0 3 96 91
0
0 0 624 270
6 74LS86
-21 -24 21 -16
4 U15D
-12 -2 16 6
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 4 11 0
1 U
3714 0 0
2
44808.6 0
0
6 74LS83
105 1247 503 0 14 29
0 2 2 2 104 114 115 116 117 113
214 102 101 100 215
0
0 0 13040 512
7 74LS83A
-24 -60 25 -52
3 U14
-10 -61 11 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 512 1 0 0 0
1 U
3406 0 0
2
44808.6 3
0
6 74LS83
105 1332 658 0 14 29
0 65 66 67 2 118 70 69 68 2
99 98 97 96 113
0
0 0 13040 512
7 74LS83A
-24 -60 25 -52
3 U16
-10 -61 11 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 0 1 0 0 0
1 U
3132 0 0
2
44808.6 2
0
7 Ground~
168 1510 754 0 1 3
0 2
0
0 0 53360 0
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3842 0 0
2
44808.6 1
0
6 74LS83
105 1429 539 0 14 29
0 104 65 66 67 2 2 2 71 2
115 116 117 118 114
0
0 0 13040 512
7 74LS83A
-24 -60 25 -52
3 U17
-10 -61 11 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 0 1 0 0 0
1 U
6183 0 0
2
44808.6 0
0
6 74LS83
105 1334 804 0 14 29
0 2 2 2 108 120 121 122 123 119
84 85 86 87 216
0
0 0 13040 512
7 74LS83A
-24 -60 25 -52
3 U13
-10 -61 11 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 512 1 0 0 0
1 U
3356 0 0
2
44808.6 0
0
6 74LS83
105 1419 959 0 14 29
0 109 110 111 2 124 105 106 107 2
92 93 94 95 119
0
0 0 13040 512
7 74LS83A
-24 -60 25 -52
3 U12
-10 -61 11 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 0 1 0 0 0
1 U
3525 0 0
2
44808.6 0
0
7 Ground~
168 1597 1157 0 1 3
0 2
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3800 0 0
2
44808.6 0
0
6 74LS83
105 1516 840 0 14 29
0 108 109 110 111 2 2 2 112 2
121 122 123 124 120
0
0 0 13040 512
7 74LS83A
-24 -60 25 -52
2 U2
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 0 1 0 0 0
1 U
346 0 0
2
44808.6 0
0
7 74LS157
122 117 742 0 14 29
0 125 217 218 2 18 2 17 219 220
2 221 16 15 222
0
0 0 13040 90
7 74LS157
-24 -60 25 -52
3 U34
53 -6 74 2
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 2 6 5 10 11 13 14
15 4 7 9 12 1 3 2 6 5
10 11 13 14 15 4 7 9 12 0
65 0 0 512 1 0 0 0
1 U
3169 0 0
2
5.89999e-315 5.26354e-315
0
10 2-In NAND~
219 1522 313 0 3 22
0 70 71 127
0
0 0 624 512
4 7400
-7 -24 21 -16
4 U35A
-11 -25 17 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 13 0
1 U
4826 0 0
2
5.89999e-315 5.30499e-315
0
5 7412~
219 1400 382 0 4 22
0 126 72 127 128
0
0 0 624 180
4 7412
-7 -24 21 -16
3 U6B
-8 -25 13 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 6 0
65 0 0 0 3 2 6 0
1 U
3971 0 0
2
5.89999e-315 5.32571e-315
0
7 Ground~
168 1303 425 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3607 0 0
2
5.89999e-315 5.34643e-315
0
7 74LS157
122 1262 334 0 14 29
0 128 223 68 224 69 225 70 226 71
2 129 130 131 132
0
0 0 13040 180
7 74LS157
-24 -60 25 -52
3 U32
-17 -61 4 -53
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 2 6 5 10 11 13 14
15 4 7 9 12 1 3 2 6 5
10 11 13 14 15 4 7 9 12 0
65 0 0 512 1 0 0 0
1 U
3506 0 0
2
5.89999e-315 5.3568e-315
0
10 Ascii Key~
169 592 253 0 11 12
0 150 151 152 153 126 154 149 155 0
0 61
0
0 0 4656 180
0
4 KBD1
32 -2 60 6
0
0
0
0
0
4 SIP8
17

0 1 2 3 4 5 6 7 8 1
2 3 4 5 6 7 8 0
0 0 0 0 1 0 0 0
3 KBD
7829 0 0
2
5.89999e-315 5.36716e-315
0
7 74LS273
150 1696 144 0 18 37
0 6 5 227 149 154 126 153 152 151
150 133 134 135 136 140 139 138 137
0
0 0 13040 782
7 74LS273
-24 -60 25 -52
3 U29
51 0 72 8
0
15 DVCC=20;GND=10;
152 %D [%20bi %10bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%20bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o] %M
0
12 type:digital
5 DIP20
37

0 1 11 18 17 14 13 8 7 4
3 19 16 15 12 9 6 5 2 1
11 18 17 14 13 8 7 4 3 19
16 15 12 9 6 5 2 0
65 0 0 512 1 0 0 0
1 U
3890 0 0
2
5.89999e-315 5.37752e-315
0
7 74LS273
150 1696 331 0 18 37
0 6 5 133 134 135 136 140 139 138
137 228 229 230 72 71 70 69 68
0
0 0 13040 782
7 74LS273
-24 -60 25 -52
3 U28
51 0 72 8
0
15 DVCC=20;GND=10;
152 %D [%20bi %10bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%20bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o] %M
0
12 type:digital
5 DIP20
37

0 1 11 18 17 14 13 8 7 4
3 19 16 15 12 9 6 5 2 1
11 18 17 14 13 8 7 4 3 19
16 15 12 9 6 5 2 0
65 0 0 512 1 0 0 0
1 U
3126 0 0
2
5.89999e-315 5.38788e-315
0
7 74LS273
150 1696 451 0 18 37
0 6 5 231 232 233 72 71 70 69
68 234 235 236 103 104 65 66 67
0
0 0 13040 782
7 74LS273
-24 -60 25 -52
3 U27
51 0 72 8
0
15 DVCC=20;GND=10;
152 %D [%20bi %10bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%20bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o] %M
0
12 type:digital
5 DIP20
37

0 1 11 18 17 14 13 8 7 4
3 19 16 15 12 9 6 5 2 1
11 18 17 14 13 8 7 4 3 19
16 15 12 9 6 5 2 0
65 0 0 512 1 0 0 0
1 U
3935 0 0
2
5.89999e-315 5.39306e-315
0
7 74LS273
150 1697 553 0 18 37
0 6 5 237 238 239 103 104 65 66
67 240 241 242 243 173 3 174 175
0
0 0 13040 782
7 74LS273
-24 -60 25 -52
3 U26
51 0 72 8
0
15 DVCC=20;GND=10;
152 %D [%20bi %10bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%20bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o] %M
0
12 type:digital
5 DIP20
37

0 1 11 18 17 14 13 8 7 4
3 19 16 15 12 9 6 5 2 1
11 18 17 14 13 8 7 4 3 19
16 15 12 9 6 5 2 0
65 0 0 512 1 0 0 0
1 U
9746 0 0
2
5.89999e-315 5.39824e-315
0
7 74LS273
150 1697 637 0 18 37
0 6 5 244 245 246 247 173 3 174
175 248 249 250 251 112 105 106 107
0
0 0 13040 782
7 74LS273
-24 -60 25 -52
3 U25
51 0 72 8
0
15 DVCC=20;GND=10;
152 %D [%20bi %10bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%20bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o] %M
0
12 type:digital
5 DIP20
37

0 1 11 18 17 14 13 8 7 4
3 19 16 15 12 9 6 5 2 1
11 18 17 14 13 8 7 4 3 19
16 15 12 9 6 5 2 0
65 0 0 512 1 0 0 0
1 U
7330 0 0
2
5.89999e-315 5.40342e-315
0
7 74LS273
150 1696 733 0 18 37
0 6 5 252 253 254 255 112 105 106
107 256 257 258 259 108 109 110 111
0
0 0 13040 782
7 74LS273
-24 -60 25 -52
3 U23
51 0 72 8
0
15 DVCC=20;GND=10;
152 %D [%20bi %10bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%20bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o] %M
0
12 type:digital
5 DIP20
37

0 1 11 18 17 14 13 8 7 4
3 19 16 15 12 9 6 5 2 1
11 18 17 14 13 8 7 4 3 19
16 15 12 9 6 5 2 0
65 0 0 512 1 0 0 0
1 U
3972 0 0
2
5.89999e-315 5.4086e-315
0
2 +V
167 321 387 0 1 3
0 6
0
0 0 54256 0
2 5V
-7 -22 7 -14
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
7818 0 0
2
5.89999e-315 5.47854e-315
0
9 CA 7-Seg~
184 111 506 0 18 19
10 260 14 14 261 262 263 13 264 172
2 2 2 2 2 2 2 2 1
0
0 0 21104 0
5 REDCA
16 -41 51 -33
5 DISP3
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
3818 0 0
2
5.89999e-315 5.47984e-315
0
6 74LS47
187 304 635 0 14 29
0 141 142 143 144 265 266 168 167 164
170 165 166 169 267
0
0 0 13040 602
6 74LS47
-21 -60 21 -52
3 U11
57 0 78 8
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
8835 0 0
2
5.89999e-315 5.48113e-315
0
9 CA 7-Seg~
184 321 508 0 18 19
10 169 166 165 170 164 167 168 268 171
2 2 2 2 2 2 2 2 1
0
0 0 21104 0
5 REDCA
16 -41 51 -33
5 DISP2
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
7484 0 0
2
5.89999e-315 5.48243e-315
0
9 CA 7-Seg~
184 541 505 0 18 19
10 161 158 157 162 156 159 160 269 163
2 2 2 2 2 2 2 2 1
0
0 0 21104 0
5 REDCA
16 -41 51 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
792 0 0
2
5.89999e-315 5.48372e-315
0
6 74LS47
187 524 637 0 14 29
0 145 146 147 148 270 271 160 159 156
162 157 158 161 272
0
0 0 13040 602
6 74LS47
-21 -60 21 -52
2 U9
60 0 74 8
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
3826 0 0
2
5.89999e-315 5.48502e-315
0
9 Inverter~
13 1617 71 0 2 22
0 155 5
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U4B
20 -8 41 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 2 4 0
1 U
7958 0 0
2
5.89999e-315 5.49408e-315
0
7 74LS157
122 549 744 0 14 29
0 125 137 26 138 25 139 24 140 23
2 148 147 146 145
0
0 0 13040 90
7 74LS157
-24 -60 25 -52
3 U30
53 -6 74 2
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 2 6 5 10 11 13 14
15 4 7 9 12 1 3 2 6 5
10 11 13 14 15 4 7 9 12 0
65 0 0 0 1 0 0 0
1 U
6736 0 0
2
5.89999e-315 5.49538e-315
0
7 74LS157
122 328 743 0 14 29
0 125 129 22 130 21 131 20 132 19
2 144 143 142 141
0
0 0 13040 90
7 74LS157
-24 -60 25 -52
3 U31
53 -6 74 2
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 2 6 5 10 11 13 14
15 4 7 9 12 1 3 2 6 5
10 11 13 14 15 4 7 9 12 0
65 0 0 0 1 0 0 0
1 U
3755 0 0
2
5.89999e-315 5.49667e-315
0
9 Resistor~
219 111 435 0 4 5
0 172 6 0 1
0
0 0 880 90
2 1k
8 0 22 8
2 R3
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
397 0 0
2
5.89999e-315 5.51286e-315
0
9 Resistor~
219 321 434 0 4 5
0 171 6 0 1
0
0 0 880 90
2 1k
8 0 22 8
2 R2
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
5190 0 0
2
5.89999e-315 5.51351e-315
0
9 Resistor~
219 541 424 0 4 5
0 163 6 0 1
0
0 0 880 90
2 1k
8 0 22 8
2 R1
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9188 0 0
2
5.89999e-315 5.51416e-315
0
368
0 1 3 0 0 8208 0 0 1 4 0 5
793 685
779 685
779 836
797 836
797 851
0 2 4 0 0 4224 0 0 1 176 0 4
827 693
827 837
815 837
815 851
1 0 2 0 0 12288 0 33 0 0 270 4
1034 759
1115 759
1115 878
1399 878
1 0 3 0 0 8320 0 20 0 0 361 3
793 707
793 595
1719 595
2 0 5 0 0 8192 0 59 0 0 332 3
1665 526
1665 494
1620 494
1 0 6 0 0 4096 0 59 0 0 242 2
1656 520
1594 520
12 4 7 0 0 8320 0 5 4 0 0 4
1139 2213
1139 2235
1186 2235
1186 2250
12 4 8 0 0 8320 0 6 7 0 0 4
1139 1964
1139 1986
1186 1986
1186 2001
12 4 9 0 0 8320 0 8 9 0 0 4
801 2173
801 2196
848 2196
848 2210
12 4 10 0 0 8320 0 11 10 0 0 4
801 1928
801 1948
848 1948
848 1965
12 4 11 0 0 8320 0 12 13 0 0 4
801 1682
801 1703
848 1703
848 1719
12 4 12 0 0 8320 0 15 14 0 0 4
801 1435
801 1458
848 1458
848 1472
6 0 2 0 0 0 0 50 0 0 14 2
121 773
121 862
4 0 2 0 0 8320 0 50 0 0 179 4
103 773
103 862
686 862
686 780
2 7 13 0 0 4224 0 2 63 0 0 2
126 607
126 542
2 0 14 0 0 4096 0 63 0 0 17 2
96 542
96 562
2 3 14 0 0 4224 0 3 63 0 0 4
96 647
96 562
102 562
102 542
1 13 15 0 0 4224 0 2 50 0 0 4
126 643
126 683
130 683
130 709
12 1 16 0 0 4224 0 50 3 0 0 4
112 709
112 690
96 690
96 683
7 0 17 0 0 8320 0 50 0 0 174 5
130 773
130 841
765 841
765 792
802 792
5 10 18 0 0 4224 0 50 4 0 0 4
112 773
112 2334
1186 2334
1186 2314
9 11 19 0 0 4224 0 70 4 0 0 4
359 774
359 2344
1195 2344
1195 2314
7 12 20 0 0 4224 0 70 4 0 0 4
341 774
341 2357
1204 2357
1204 2314
5 13 21 0 0 4224 0 70 4 0 0 4
323 774
323 2368
1213 2368
1213 2314
10 3 22 0 0 12416 0 9 70 0 0 4
848 2274
848 2292
305 2292
305 774
9 11 23 0 0 4224 0 69 9 0 0 4
580 775
580 2304
857 2304
857 2274
12 7 24 0 0 12416 0 9 69 0 0 4
866 2274
866 2313
562 2313
562 775
13 5 25 0 0 12416 0 9 69 0 0 4
875 2274
875 2323
544 2323
544 775
13 3 26 0 0 8320 0 32 69 0 0 4
1062 1178
1062 1297
526 1297
526 775
10 8 27 0 0 16512 0 10 4 0 0 6
848 2029
848 2049
990 2049
990 2079
1222 2079
1222 2250
10 0 28 0 0 12288 0 5 0 0 48 4
1103 2213
1103 2231
1047 2231
1047 1978
2 0 2 0 0 0 0 4 0 0 33 2
1168 2250
1168 2223
1 0 2 0 0 0 0 4 0 0 39 3
1159 2250
1159 2223
1240 2223
3 0 7 0 0 0 0 4 0 0 7 2
1177 2250
1177 2235
8 0 27 0 0 0 0 5 0 0 30 3
1157 2149
1157 2148
1222 2148
7 0 29 0 0 8192 0 5 0 0 40 3
1148 2149
1148 2135
1213 2135
6 0 30 0 0 8192 0 5 0 0 41 3
1139 2149
1139 2125
1204 2125
5 0 31 0 0 8192 0 5 0 0 42 3
1130 2149
1130 2114
1195 2114
9 0 2 0 0 0 0 4 0 0 59 4
1240 2250
1240 2102
1026 2102
1026 1820
13 7 29 0 0 4224 0 7 4 0 0 2
1213 2065
1213 2250
12 6 30 0 0 4224 0 7 4 0 0 2
1204 2065
1204 2250
11 5 31 0 0 4224 0 7 4 0 0 2
1195 2065
1195 2250
4 0 2 0 0 0 0 5 0 0 45 3
1121 2149
1121 2119
1094 2119
3 0 2 0 0 0 0 5 0 0 45 3
1112 2149
1112 2128
1094 2128
1 0 2 0 0 0 0 5 0 0 39 2
1094 2149
1094 2102
2 0 28 0 0 0 0 5 0 0 31 3
1103 2149
1103 2138
1047 2138
10 8 32 0 0 8320 0 13 7 0 0 4
848 1783
848 1800
1222 1800
1222 2001
0 10 28 0 0 8320 0 0 6 110 0 5
708 1559
1047 1559
1047 1978
1103 1978
1103 1964
9 0 2 0 0 0 0 7 0 0 99 5
1240 2001
1240 1852
1026 1852
1026 1607
902 1607
2 0 2 0 0 0 0 7 0 0 51 2
1168 2001
1168 1973
1 0 2 0 0 0 0 7 0 0 49 3
1159 2001
1159 1973
1240 1973
3 0 8 0 0 0 0 7 0 0 8 2
1177 2001
1177 1986
8 0 32 0 0 0 0 6 0 0 47 3
1157 1900
1157 1896
1222 1896
7 0 33 0 0 8192 0 6 0 0 57 3
1148 1900
1148 1886
1213 1886
6 0 34 0 0 8192 0 6 0 0 58 3
1139 1900
1139 1876
1204 1876
5 0 2 0 0 0 0 6 0 0 59 3
1130 1900
1130 1865
1195 1865
10 7 33 0 0 12416 0 14 7 0 0 4
848 1536
848 1550
1213 1550
1213 2001
10 6 34 0 0 12416 0 19 7 0 0 4
848 1287
848 1308
1204 1308
1204 2001
0 5 2 0 0 0 0 0 7 49 0 3
1026 1820
1195 1820
1195 2001
4 0 2 0 0 0 0 6 0 0 62 3
1121 1900
1121 1870
1094 1870
3 0 2 0 0 0 0 6 0 0 62 3
1112 1900
1112 1879
1094 1879
1 0 2 0 0 0 0 6 0 0 49 2
1094 1900
1094 1852
2 0 28 0 0 0 0 6 0 0 48 3
1103 1900
1103 1890
1047 1890
12 8 35 0 0 12416 0 32 9 0 0 6
1053 1178
1053 1215
953 1215
953 2074
884 2074
884 2210
9 0 2 0 0 0 0 9 0 0 82 4
902 2210
902 2061
688 2061
688 1816
2 0 2 0 0 0 0 9 0 0 67 2
830 2210
830 2182
1 0 2 0 0 0 0 9 0 0 65 3
821 2210
821 2182
902 2182
3 0 9 0 0 0 0 9 0 0 9 2
839 2210
839 2196
8 0 35 0 0 0 0 8 0 0 64 3
819 2109
819 2101
884 2101
7 0 36 0 0 8192 0 8 0 0 73 3
810 2109
810 2095
875 2095
6 0 37 0 0 8192 0 8 0 0 74 3
801 2109
801 2085
866 2085
5 0 38 0 0 8192 0 8 0 0 75 3
792 2109
792 2074
857 2074
13 7 36 0 0 4224 0 10 9 0 0 2
875 2029
875 2210
12 6 37 0 0 4224 0 10 9 0 0 2
866 2029
866 2210
11 5 38 0 0 4224 0 10 9 0 0 2
857 2029
857 2210
10 0 28 0 0 0 0 8 0 0 93 4
765 2173
765 2191
708 2191
708 1946
4 0 2 0 0 0 0 8 0 0 79 3
783 2109
783 2079
756 2079
3 0 2 0 0 0 0 8 0 0 79 3
774 2109
774 2088
756 2088
1 0 2 0 0 0 0 8 0 0 65 2
756 2109
756 2061
2 0 28 0 0 0 0 8 0 0 76 3
765 2109
765 2098
708 2098
11 8 39 0 0 12416 0 32 10 0 0 6
1044 1178
1044 1207
945 1207
945 1828
884 1828
884 1965
9 0 2 0 0 0 0 10 0 0 99 4
902 1965
902 1816
688 1816
688 1570
2 0 2 0 0 0 0 10 0 0 84 2
830 1965
830 1937
1 0 2 0 0 0 0 10 0 0 82 3
821 1965
821 1937
902 1937
3 0 10 0 0 0 0 10 0 0 10 2
839 1965
839 1948
8 0 39 0 0 0 0 11 0 0 81 3
819 1864
819 1856
884 1856
7 0 40 0 0 8192 0 11 0 0 90 3
810 1864
810 1850
875 1850
6 0 41 0 0 8192 0 11 0 0 91 3
801 1864
801 1840
866 1840
5 0 42 0 0 8192 0 11 0 0 92 3
792 1864
792 1829
857 1829
13 7 40 0 0 4224 0 13 10 0 0 2
875 1783
875 1965
12 6 41 0 0 4224 0 13 10 0 0 2
866 1783
866 1965
11 5 42 0 0 4224 0 13 10 0 0 2
857 1783
857 1965
10 0 28 0 0 0 0 11 0 0 110 4
765 1928
765 1946
708 1946
708 1700
4 0 2 0 0 0 0 11 0 0 96 3
783 1864
783 1834
756 1834
3 0 2 0 0 0 0 11 0 0 96 3
774 1864
774 1843
756 1843
1 0 2 0 0 0 0 11 0 0 82 2
756 1864
756 1816
2 0 28 0 0 0 0 11 0 0 93 3
765 1864
765 1853
708 1853
8 10 43 0 0 12416 0 13 32 0 0 6
884 1719
884 1582
937 1582
937 1199
1035 1199
1035 1178
9 0 2 0 0 0 0 13 0 0 122 4
902 1719
902 1570
688 1570
688 1324
2 0 2 0 0 0 0 13 0 0 101 2
830 1719
830 1691
1 0 2 0 0 0 0 13 0 0 99 3
821 1719
821 1691
902 1691
3 0 11 0 0 0 0 13 0 0 11 2
839 1719
839 1703
8 0 43 0 0 0 0 12 0 0 98 3
819 1618
819 1613
884 1613
7 0 44 0 0 8192 0 12 0 0 107 3
810 1618
810 1604
875 1604
6 0 45 0 0 8192 0 12 0 0 108 3
801 1618
801 1594
866 1594
5 0 46 0 0 8192 0 12 0 0 109 3
792 1618
792 1583
857 1583
13 7 44 0 0 4224 0 14 13 0 0 2
875 1536
875 1719
12 6 45 0 0 4224 0 14 13 0 0 2
866 1536
866 1719
11 5 46 0 0 4224 0 14 13 0 0 2
857 1536
857 1719
10 0 28 0 0 0 0 12 0 0 128 4
765 1682
765 1700
708 1700
708 1453
4 0 2 0 0 0 0 12 0 0 113 3
783 1618
783 1588
756 1588
3 0 2 0 0 0 0 12 0 0 113 3
774 1618
774 1597
756 1597
1 0 2 0 0 0 0 12 0 0 99 2
756 1618
756 1570
2 0 28 0 0 0 0 12 0 0 110 3
765 1618
765 1607
708 1607
2 0 2 0 0 0 0 14 0 0 116 2
830 1472
830 1445
1 0 2 0 0 0 0 14 0 0 122 3
821 1472
821 1445
902 1445
3 0 12 0 0 0 0 14 0 0 12 2
839 1472
839 1458
8 0 47 0 0 8192 0 15 0 0 124 3
819 1371
819 1366
884 1366
7 0 48 0 0 8192 0 15 0 0 125 3
810 1371
810 1357
875 1357
6 0 49 0 0 8192 0 15 0 0 126 3
801 1371
801 1347
866 1347
5 0 50 0 0 8192 0 15 0 0 127 3
792 1371
792 1336
857 1336
9 0 2 0 0 0 0 14 0 0 140 5
902 1472
902 1324
688 1324
688 1044
752 1044
9 0 2 0 0 0 0 19 0 0 136 3
902 1223
902 1204
857 1204
13 8 47 0 0 12416 0 24 14 0 0 6
893 1108
893 1199
927 1199
927 1338
884 1338
884 1472
13 7 48 0 0 4224 0 19 14 0 0 2
875 1287
875 1472
12 6 49 0 0 4224 0 19 14 0 0 2
866 1287
866 1472
11 5 50 0 0 4224 0 19 14 0 0 2
857 1287
857 1472
10 1 28 0 0 0 0 15 0 0 137 4
765 1435
765 1453
708 1453
708 1212
4 0 2 0 0 0 0 15 0 0 131 3
783 1371
783 1341
756 1341
3 0 2 0 0 0 0 15 0 0 131 3
774 1371
774 1350
756 1350
1 0 2 0 0 0 0 15 0 0 122 2
756 1371
756 1324
2 0 28 0 0 0 0 15 0 0 128 3
765 1371
765 1360
708 1360
3 0 51 0 0 4096 0 19 0 0 134 2
839 1223
839 1213
12 4 51 0 0 8320 0 18 19 0 0 4
801 1194
801 1213
848 1213
848 1223
2 0 2 0 0 0 0 19 0 0 136 2
830 1223
830 1204
1 0 2 0 0 0 0 19 0 0 142 3
821 1223
821 1204
857 1204
10 1 28 0 0 0 0 18 16 0 0 4
765 1194
765 1212
708 1212
708 970
4 0 2 0 0 0 0 18 0 0 140 3
783 1130
783 1100
752 1100
3 0 2 0 0 0 0 18 0 0 140 3
774 1130
774 1109
752 1109
1 0 2 0 0 0 0 18 0 0 153 3
756 1130
752 1130
752 1028
2 0 28 0 0 0 0 18 0 0 137 3
765 1130
765 1119
708 1119
5 0 2 0 0 0 0 19 0 0 143 5
857 1223
857 1133
843 1133
843 1106
792 1106
5 0 2 0 0 0 0 18 0 0 153 2
792 1130
792 1028
6 0 52 0 0 8192 0 18 0 0 147 3
801 1130
801 1113
866 1113
7 0 53 0 0 8192 0 18 0 0 148 3
810 1130
810 1118
875 1118
8 0 54 0 0 8192 0 18 0 0 149 3
819 1130
819 1124
884 1124
10 6 52 0 0 4224 0 24 19 0 0 2
866 1108
866 1223
11 7 53 0 0 4224 0 24 19 0 0 2
875 1108
875 1223
12 8 54 0 0 4224 0 24 19 0 0 2
884 1108
884 1223
3 0 2 0 0 0 0 24 0 0 153 2
857 1044
857 1028
2 0 2 0 0 0 0 24 0 0 153 2
848 1044
848 1028
1 0 2 0 0 0 0 24 0 0 153 2
839 1044
839 1028
4 1 2 0 0 0 0 24 17 0 0 4
866 1044
866 1028
752 1028
752 952
3 5 55 0 0 4224 0 1 24 0 0 4
806 903
806 1018
875 1018
875 1044
3 6 56 0 0 4224 0 30 24 0 0 4
853 883
853 1009
884 1009
884 1044
3 7 57 0 0 4224 0 31 24 0 0 4
896 884
896 1010
893 1010
893 1044
3 8 58 0 0 4224 0 29 24 0 0 4
938 884
938 1020
902 1020
902 1044
9 14 59 0 0 12416 0 24 32 0 0 5
920 1044
942 1044
942 1188
1089 1188
1089 1178
8 0 2 0 0 0 0 32 0 0 162 2
1071 1114
1071 1077
7 0 2 0 0 0 0 32 0 0 162 2
1062 1114
1062 1077
6 0 2 0 0 0 0 32 0 0 162 2
1053 1114
1053 1077
5 0 2 0 0 0 0 32 0 0 285 3
1044 1114
1044 1077
1597 1077
4 3 60 0 0 8320 0 32 28 0 0 4
1035 1114
1035 1098
1118 1098
1118 1059
3 3 61 0 0 8320 0 32 25 0 0 4
1026 1114
1026 1087
1076 1087
1076 1059
2 3 62 0 0 4224 0 32 27 0 0 4
1017 1114
1017 1082
1033 1082
1033 1058
1 3 63 0 0 4224 0 32 26 0 0 4
1008 1114
1008 1082
991 1082
991 1057
0 9 17 0 0 0 0 0 32 171 0 4
956 999
956 1093
1089 1093
1089 1114
2 0 17 0 0 0 0 25 0 0 171 2
1067 1010
1067 999
2 0 17 0 0 0 0 27 0 0 171 2
1024 1009
1024 999
2 0 17 0 0 0 0 26 0 0 171 2
982 1008
982 999
0 2 17 0 0 128 0 0 28 174 0 4
914 817
914 999
1109 999
1109 1010
2 0 17 0 0 0 0 31 0 0 174 2
887 835
887 817
2 0 17 0 0 0 0 30 0 0 174 2
844 834
844 817
3 2 17 0 0 0 0 20 29 0 0 4
802 752
802 817
929 817
929 835
1 10 64 0 0 8320 0 23 33 0 0 4
901 693
922 693
922 786
970 786
2 2 4 0 0 128 0 23 20 0 0 3
865 693
811 693
811 707
10 10 2 0 0 0 0 50 70 0 0 3
157 779
157 780
368 780
10 0 2 0 0 0 0 69 0 0 179 2
589 781
589 780
10 1 2 0 0 128 0 70 21 0 0 3
368 780
686 780
686 766
1 0 65 0 0 4096 0 43 0 0 236 3
1364 622
1529 622
1529 507
2 0 66 0 0 4096 0 43 0 0 235 3
1364 631
1535 631
1535 510
3 0 67 0 0 4096 0 43 0 0 234 3
1364 640
1542 640
1542 513
2 0 5 0 0 4096 0 58 0 0 332 3
1664 424
1664 371
1620 371
10 18 68 0 0 4096 0 58 57 0 0 2
1736 424
1736 368
9 17 69 0 0 4096 0 58 57 0 0 2
1727 424
1727 368
8 16 70 0 0 4096 0 58 57 0 0 2
1718 424
1718 368
7 15 71 0 0 4096 0 58 57 0 0 2
1709 424
1709 368
6 14 72 0 0 4096 0 58 57 0 0 2
1700 424
1700 368
1 11 73 0 0 8320 0 30 33 0 0 3
862 834
862 795
970 795
12 1 74 0 0 4224 0 33 31 0 0 3
970 804
905 804
905 835
13 1 75 0 0 4224 0 33 29 0 0 3
970 813
947 813
947 835
10 1 76 0 0 4224 0 34 26 0 0 3
1138 941
1000 941
1000 1008
11 1 77 0 0 4224 0 34 27 0 0 3
1138 950
1042 950
1042 1009
12 1 78 0 0 4224 0 34 25 0 0 3
1138 959
1085 959
1085 1010
13 1 79 0 0 8320 0 34 28 0 0 3
1138 968
1127 968
1127 1010
2 3 80 0 0 8320 0 33 36 0 0 5
1034 768
1059 768
1059 686
994 686
994 670
3 3 81 0 0 8320 0 33 37 0 0 5
1034 777
1069 777
1069 676
1037 676
1037 671
3 4 82 0 0 4224 0 35 33 0 0 3
1079 671
1079 786
1034 786
9 14 83 0 0 8320 0 33 34 0 0 4
1034 840
1103 840
1103 995
1138 995
5 10 84 0 0 4224 0 33 46 0 0 2
1034 795
1302 795
6 11 85 0 0 4224 0 33 46 0 0 2
1034 804
1302 804
7 12 86 0 0 4224 0 33 46 0 0 2
1034 813
1302 813
8 13 87 0 0 4224 0 33 46 0 0 2
1034 822
1302 822
1 3 88 0 0 8320 0 34 40 0 0 5
1202 914
1228 914
1228 768
1130 768
1130 739
2 3 89 0 0 8320 0 34 39 0 0 5
1202 923
1240 923
1240 759
1172 759
1172 740
3 3 90 0 0 8320 0 34 38 0 0 5
1202 932
1249 932
1249 750
1215 750
1215 741
4 3 91 0 0 8320 0 34 41 0 0 3
1202 941
1257 941
1257 741
9 0 3 0 0 0 0 34 0 0 4 3
1202 995
1278 995
1278 595
5 10 92 0 0 4224 0 34 47 0 0 2
1202 950
1387 950
6 11 93 0 0 4224 0 34 47 0 0 2
1202 959
1387 959
12 7 94 0 0 4224 0 47 34 0 0 2
1387 968
1202 968
13 8 95 0 0 4224 0 47 34 0 0 2
1387 977
1202 977
2 13 96 0 0 8320 0 41 43 0 0 3
1248 692
1248 676
1300 676
2 12 97 0 0 8320 0 38 43 0 0 3
1206 692
1206 667
1300 667
2 11 98 0 0 8320 0 39 43 0 0 3
1163 691
1163 658
1300 658
2 10 99 0 0 8320 0 40 43 0 0 3
1121 690
1121 649
1300 649
2 13 100 0 0 8320 0 35 42 0 0 3
1070 622
1070 521
1215 521
2 12 101 0 0 8320 0 37 42 0 0 3
1028 622
1028 512
1215 512
2 11 102 0 0 8320 0 36 42 0 0 3
985 621
985 503
1215 503
1 0 3 0 0 0 0 41 0 0 4 2
1266 692
1266 595
1 0 3 0 0 0 0 38 0 0 4 2
1224 692
1224 595
1 0 3 0 0 0 0 39 0 0 4 2
1181 691
1181 595
1 0 3 0 0 0 0 40 0 0 4 2
1139 690
1139 595
1 0 3 0 0 0 0 35 0 0 4 2
1088 622
1088 595
1 0 3 0 0 0 0 37 0 0 4 2
1046 622
1046 595
1 0 3 0 0 0 0 36 0 0 4 2
1003 621
1003 595
2 0 72 0 0 4224 0 52 0 0 188 2
1424 382
1700 382
14 6 103 0 0 12416 0 58 59 0 0 4
1700 488
1700 503
1701 503
1701 526
0 4 104 0 0 8192 0 0 42 237 0 5
1476 503
1476 481
1346 481
1346 494
1279 494
6 0 70 0 0 8320 0 43 0 0 292 3
1364 667
1550 667
1550 399
7 0 69 0 0 8192 0 43 0 0 291 3
1364 676
1557 676
1557 405
8 0 68 0 0 8192 0 43 0 0 243 3
1364 685
1562 685
1562 411
8 0 71 0 0 8192 0 45 0 0 293 3
1461 566
1500 566
1500 394
4 0 67 0 0 12416 0 45 0 0 367 4
1461 530
1494 530
1494 513
1736 513
3 0 66 0 0 12416 0 45 0 0 364 4
1461 521
1487 521
1487 510
1727 510
2 0 65 0 0 12416 0 45 0 0 363 4
1461 512
1481 512
1481 507
1718 507
1 0 104 0 0 4224 0 45 0 0 362 2
1461 503
1709 503
2 0 71 0 0 0 0 51 0 0 293 2
1548 322
1548 394
1 0 70 0 0 0 0 51 0 0 292 3
1548 304
1557 304
1557 399
1 0 6 0 0 0 0 58 0 0 242 4
1655 418
1609 418
1609 426
1594 426
1 0 6 0 0 0 0 60 0 0 242 2
1656 604
1594 604
1 0 6 0 0 8192 0 61 0 0 319 3
1655 700
1594 700
1594 225
3 0 68 0 0 12416 0 54 0 0 184 4
1288 356
1348 356
1348 411
1736 411
6 0 105 0 0 4224 0 47 0 0 357 4
1451 968
1770 968
1770 693
1718 693
7 0 106 0 0 4224 0 47 0 0 356 4
1451 977
1777 977
1777 686
1727 686
8 0 107 0 0 4224 0 47 0 0 365 4
1451 986
1786 986
1786 679
1736 679
1 0 108 0 0 8192 0 49 0 0 271 3
1548 804
1558 804
1558 779
2 0 109 0 0 4096 0 49 0 0 276 2
1548 813
1718 813
3 0 110 0 0 4096 0 49 0 0 277 2
1548 822
1727 822
4 0 111 0 0 4096 0 49 0 0 278 2
1548 831
1736 831
8 0 112 0 0 8320 0 49 0 0 358 4
1548 867
1576 867
1576 694
1709 694
14 9 113 0 0 8320 0 43 42 0 0 4
1300 703
1287 703
1287 548
1279 548
3 0 2 0 0 0 0 42 0 0 255 2
1279 485
1312 485
2 0 2 0 0 0 0 42 0 0 255 2
1279 476
1312 476
1 0 2 0 0 0 0 42 0 0 266 4
1279 467
1312 467
1312 600
1510 600
14 5 114 0 0 4224 0 45 42 0 0 4
1397 584
1297 584
1297 503
1279 503
10 6 115 0 0 12416 0 45 42 0 0 4
1397 530
1383 530
1383 512
1279 512
11 7 116 0 0 12416 0 45 42 0 0 4
1397 539
1377 539
1377 521
1279 521
12 8 117 0 0 12416 0 45 42 0 0 4
1397 548
1370 548
1370 530
1279 530
9 0 2 0 0 0 0 43 0 0 266 2
1364 703
1510 703
4 0 2 0 0 0 0 43 0 0 266 2
1364 649
1510 649
13 5 118 0 0 8320 0 45 43 0 0 4
1397 557
1386 557
1386 658
1364 658
6 0 2 0 0 0 0 45 0 0 266 2
1461 548
1510 548
7 0 2 0 0 0 0 45 0 0 266 2
1461 557
1510 557
9 0 2 0 0 0 0 45 0 0 266 2
1461 584
1510 584
5 1 2 0 0 128 0 45 44 0 0 3
1461 539
1510 539
1510 748
14 9 119 0 0 8320 0 47 46 0 0 4
1387 1004
1374 1004
1374 849
1366 849
3 0 2 0 0 0 0 46 0 0 270 2
1366 786
1399 786
2 0 2 0 0 0 0 46 0 0 270 2
1366 777
1399 777
1 0 2 0 0 0 0 46 0 0 285 4
1366 768
1399 768
1399 901
1597 901
4 15 108 0 0 12416 0 46 61 0 0 5
1366 795
1410 795
1410 779
1709 779
1709 770
14 5 120 0 0 4224 0 49 46 0 0 4
1484 885
1384 885
1384 804
1366 804
10 6 121 0 0 12416 0 49 46 0 0 4
1484 831
1470 831
1470 813
1366 813
11 7 122 0 0 12416 0 49 46 0 0 4
1484 840
1464 840
1464 822
1366 822
12 8 123 0 0 12416 0 49 46 0 0 4
1484 849
1457 849
1457 831
1366 831
1 16 109 0 0 4224 0 47 61 0 0 3
1451 923
1718 923
1718 770
2 17 110 0 0 4224 0 47 61 0 0 3
1451 932
1727 932
1727 770
3 18 111 0 0 4224 0 47 61 0 0 3
1451 941
1736 941
1736 770
9 0 2 0 0 0 0 47 0 0 285 2
1451 1004
1597 1004
4 0 2 0 0 0 0 47 0 0 285 2
1451 950
1597 950
13 5 124 0 0 8320 0 49 47 0 0 4
1484 858
1473 858
1473 959
1451 959
6 0 2 0 0 0 0 49 0 0 285 2
1548 849
1597 849
7 0 2 0 0 0 0 49 0 0 285 2
1548 858
1597 858
9 0 2 0 0 0 0 49 0 0 285 2
1548 885
1597 885
5 1 2 0 0 0 0 49 48 0 0 3
1548 840
1597 840
1597 1151
0 1 125 0 0 4096 0 0 50 307 0 3
287 802
76 802
76 773
1 0 126 0 0 8192 0 52 0 0 288 3
1424 391
1573 391
1573 189
1 0 126 0 0 0 0 22 0 0 326 3
1431 190
1573 190
1573 98
3 3 127 0 0 4224 0 51 52 0 0 4
1497 313
1431 313
1431 373
1424 373
4 1 128 0 0 8320 0 52 54 0 0 3
1373 382
1373 374
1288 374
5 0 69 0 0 12416 0 54 0 0 185 4
1288 338
1444 338
1444 405
1727 405
7 0 70 0 0 0 0 54 0 0 186 4
1288 320
1451 320
1451 399
1718 399
9 0 71 0 0 12416 0 54 0 0 187 4
1288 302
1459 302
1459 394
1709 394
11 2 129 0 0 4224 0 54 70 0 0 5
1224 356
451 356
451 825
296 825
296 774
12 4 130 0 0 4224 0 54 70 0 0 5
1224 338
437 338
437 813
314 813
314 774
13 6 131 0 0 4224 0 54 70 0 0 5
1224 320
422 320
422 790
332 790
332 774
14 8 132 0 0 4224 0 54 70 0 0 5
1224 302
407 302
407 785
350 785
350 774
3 11 133 0 0 4224 0 57 56 0 0 2
1673 304
1673 181
4 12 134 0 0 4224 0 57 56 0 0 2
1682 304
1682 181
5 13 135 0 0 4224 0 57 56 0 0 2
1691 304
1691 181
6 14 136 0 0 4224 0 57 56 0 0 2
1700 304
1700 181
10 1 2 0 0 0 0 54 53 0 0 3
1294 293
1303 293
1303 419
0 2 137 0 0 12416 0 0 69 368 0 7
1736 220
1495 220
1495 272
667 272
667 809
517 809
517 775
0 4 138 0 0 12416 0 0 69 355 0 7
1727 213
1480 213
1480 262
657 262
657 797
535 797
535 775
0 6 139 0 0 8320 0 0 69 310 0 6
1473 207
1473 250
650 250
650 791
553 791
553 775
0 8 140 0 0 8320 0 0 69 309 0 6
1463 198
1463 239
638 239
638 786
571 786
571 775
0 1 125 0 0 4096 0 0 70 308 0 3
510 802
287 802
287 774
4 1 125 0 0 4224 0 22 69 0 0 7
1380 199
859 199
859 414
661 414
661 802
508 802
508 775
2 0 140 0 0 0 0 22 0 0 353 4
1431 199
1463 199
1463 198
1709 198
3 0 139 0 0 0 0 22 0 0 354 4
1431 208
1473 208
1473 207
1718 207
14 1 141 0 0 4224 0 70 64 0 0 4
359 710
359 680
345 680
345 672
13 2 142 0 0 4224 0 70 64 0 0 4
341 710
341 680
336 680
336 672
12 3 143 0 0 4224 0 70 64 0 0 4
323 710
323 680
327 680
327 672
11 4 144 0 0 4224 0 70 64 0 0 4
305 710
305 680
318 680
318 672
14 1 145 0 0 4224 0 69 67 0 0 4
580 711
580 682
565 682
565 674
13 2 146 0 0 4224 0 69 67 0 0 4
562 711
562 682
556 682
556 674
12 3 147 0 0 4224 0 69 67 0 0 4
544 711
544 682
547 682
547 674
11 4 148 0 0 4224 0 69 67 0 0 4
526 711
526 682
538 682
538 674
0 1 6 0 0 0 0 0 56 320 0 3
1594 225
1594 111
1655 111
1 1 6 0 0 4224 0 62 57 0 0 5
321 396
1317 396
1317 225
1655 225
1655 298
7 4 149 0 0 8320 0 55 56 0 0 4
605 229
605 93
1682 93
1682 117
1 10 150 0 0 8320 0 55 56 0 0 4
569 229
569 93
1736 93
1736 117
2 9 151 0 0 8320 0 55 56 0 0 4
575 229
575 93
1727 93
1727 117
3 8 152 0 0 8320 0 55 56 0 0 4
581 229
581 93
1718 93
1718 117
4 7 153 0 0 8320 0 55 56 0 0 4
587 229
587 93
1709 93
1709 117
5 6 126 0 0 8320 0 55 56 0 0 4
593 229
593 98
1700 98
1700 117
6 5 154 0 0 8320 0 55 56 0 0 4
599 229
599 103
1691 103
1691 117
8 1 155 0 0 8320 0 55 68 0 0 4
611 229
611 51
1620 51
1620 53
2 0 5 0 0 0 0 60 0 0 332 3
1665 610
1665 588
1620 588
2 0 5 0 0 4096 0 57 0 0 332 3
1664 304
1664 196
1620 196
2 2 5 0 0 0 0 56 68 0 0 4
1664 117
1664 106
1620 106
1620 89
2 2 5 0 0 12416 0 61 68 0 0 4
1664 706
1664 687
1620 687
1620 89
2 1 6 0 0 0 0 73 62 0 0 3
541 406
541 396
321 396
9 5 156 0 0 12416 0 67 66 0 0 4
547 604
547 577
544 577
544 541
11 3 157 0 0 12416 0 67 66 0 0 4
529 604
529 577
532 577
532 541
12 2 158 0 0 4224 0 67 66 0 0 4
520 604
520 565
526 565
526 541
8 6 159 0 0 4224 0 67 66 0 0 4
556 604
556 565
550 565
550 541
7 7 160 0 0 4224 0 67 66 0 0 4
565 604
565 555
556 555
556 541
13 1 161 0 0 4224 0 67 66 0 0 4
511 604
511 555
520 555
520 541
10 4 162 0 0 4224 0 67 66 0 0 2
538 604
538 541
9 1 163 0 0 4224 0 66 73 0 0 2
541 469
541 442
2 1 6 0 0 0 0 71 62 0 0 3
111 417
111 396
321 396
2 1 6 0 0 0 0 72 62 0 0 2
321 416
321 396
9 5 164 0 0 4224 0 64 65 0 0 4
327 602
327 571
324 571
324 544
11 3 165 0 0 4224 0 64 65 0 0 4
309 602
309 571
312 571
312 544
12 2 166 0 0 4224 0 64 65 0 0 4
300 602
300 559
306 559
306 544
8 6 167 0 0 4224 0 64 65 0 0 4
336 602
336 559
330 559
330 544
7 7 168 0 0 4224 0 64 65 0 0 4
345 602
345 549
336 549
336 544
13 1 169 0 0 4224 0 64 65 0 0 4
291 602
291 549
300 549
300 544
10 4 170 0 0 4224 0 64 65 0 0 2
318 602
318 544
9 1 171 0 0 4224 0 65 72 0 0 2
321 472
321 452
9 1 172 0 0 4224 0 63 71 0 0 2
111 470
111 453
7 15 140 0 0 0 0 57 56 0 0 2
1709 304
1709 181
8 16 139 0 0 0 0 57 56 0 0 2
1718 304
1718 181
9 17 138 0 0 0 0 57 56 0 0 2
1727 304
1727 181
17 9 106 0 0 0 0 60 61 0 0 4
1728 674
1728 686
1727 686
1727 706
16 8 105 0 0 0 0 60 61 0 0 4
1719 674
1719 693
1718 693
1718 706
7 15 112 0 0 0 0 61 60 0 0 4
1709 706
1709 694
1710 694
1710 674
15 7 173 0 0 4224 0 59 60 0 0 2
1710 590
1710 610
17 9 174 0 0 4224 0 59 60 0 0 2
1728 590
1728 610
16 8 3 0 0 0 0 59 60 0 0 6
1719 590
1719 595
1718 595
1718 595
1719 595
1719 610
15 7 104 0 0 0 0 58 59 0 0 4
1709 488
1709 503
1710 503
1710 526
16 8 65 0 0 0 0 58 59 0 0 4
1718 488
1718 507
1719 507
1719 526
17 9 66 0 0 0 0 58 59 0 0 4
1727 488
1727 510
1728 510
1728 526
10 18 107 0 0 0 0 61 60 0 0 4
1736 706
1736 679
1737 679
1737 674
10 18 175 0 0 4224 0 60 59 0 0 2
1737 610
1737 590
10 18 67 0 0 0 0 59 58 0 0 4
1737 526
1737 513
1736 513
1736 488
18 10 137 0 0 0 0 56 57 0 0 2
1736 181
1736 304
20
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 50
577 838 798 902
587 846 787 894
50 When op is neg -> C7 is 0
otherwise, C7 is itself
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 15
53 575 194 599
63 583 183 599
15 displays 1 or -
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 134
1254 1977 1459 2121
1264 1985 1448 2097
134 This s4 is 2nd
least significant digit
in hundredth place
i.e, if ON - hundredth 
place is >=2 but here
max hundredth place is
1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 67
673 616 934 680
683 624 923 672
67 select line to do 2s comp of C
1 when op is - & C7 is 0
res is <0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 13
703 991 828 1015
713 999 817 1015
13 resh - Binary
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 13
1110 1096 1235 1120
1120 1104 1224 1120
13 resl - Binary
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
945 740 982 764
955 748 971 764
2 Ch
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1111 901 1148 925
1121 909 1137 925
2 Cl
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 36
1161 1004 1350 1048
1171 1012 1339 1044
36 Add 1 incase of - for
2s complement
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 41
1090 597 1279 641
1100 605 1268 637
41 2s complement of B
incase of - operation
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 44
354 676 567 720
364 684 556 716
44 MUX to current number or
res when pressed =
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 17
1222 168 1379 192
1232 176 1368 192
17 Logic to detect =
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 57
1007 299 1212 363
1017 307 1201 355
57 MUX to 15 or previous 
number if previous is a 
number
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1366 922 1403 946
1376 930 1392 946
2 Al
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1281 764 1318 788
1291 772 1307 788
2 Ah
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1279 615 1316 639
1289 623 1305 639
2 Bl
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1189 462 1226 486
1199 470 1215 486
2 Bh
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 16
981 568 1130 592
991 576 1119 592
16 +/- Sign 1 for -
-37 0 0 0 700 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 23
37 86 574 149
52 94 558 135
23 Double Digit Calculator
-37 0 0 0 700 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 23
37 87 574 150
52 95 558 136
23 _______________________
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
